module processor_core
    (
        input wire clk,rst
    );

endmodule
