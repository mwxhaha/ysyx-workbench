module my_not(a,b);
  input  a;
  output b;

  assign b = ~a;
endmodule
