`include "config.vh"
`include "inst.vh"

module exu_mem (
    input wire clk,
    input wire rst,
    input wire [`INST_NUM_WIDTH-1:0] inst_num,
    input wire [`INST_TYPE_WIDTH-1:0] inst_type,
    input wire [`IMM_WIDTH-1:0] imm,
    input wire [`ISA_WIDTH-1:0] pc_out,
    input wire [`ISA_WIDTH-1:0] src1,
    input wire [`ISA_WIDTH-1:0] src2,
    input wire [`ISA_WIDTH-1:0] mem_r,
    output wire [`ISA_WIDTH-1:0] mem_w,
    output wire [`ISA_WIDTH-1:0] mem_addr,
    output wire [`MEM_MASK_WIDTH-1:0] mem_mask,
    output wire mem_r_en,
    output wire mem_w_en,
    input wire [`ISA_WIDTH-1:0] alu_result
);

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(`ISA_WIDTH)
    ) muxkeywithdefault_mem_w (
        .out(mem_w),
        .key(inst_num),
        .default_out(`ISA_WIDTH'b0),
        .lut({
            `INST_NUM_WIDTH'd`lui,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`auipc,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`jal,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`jalr,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`beq,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`bne,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`blt,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`bge,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`bltu,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`bgeu,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`lb,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`lh,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`lw,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`lbu,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`lhu,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`sb,
            {{`ISA_WIDTH - 8{1'b0}}, src2[7:0]},
            `INST_NUM_WIDTH'd`sh,
            {{`ISA_WIDTH - 16{1'b0}}, src2[15:0]},
            `INST_NUM_WIDTH'd`sw,
            {{`ISA_WIDTH - 32{1'b0}}, src2[31:0]},
            `INST_NUM_WIDTH'd`addi,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`slti,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`sltiu,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`xori,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`ori,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`andi,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`slli,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`srli,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`srai,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`add,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`sub,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`sll,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`slt,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`sltu,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`ixor,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`srl,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`sra,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`ior,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`iand,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`ebreak,
            `ISA_WIDTH'b0
        })
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(`ISA_WIDTH)
    ) muxkeywithdefault_mem_addr (
        .out(mem_addr),
        .key(inst_num),
        .default_out(`BASE_ADDR),
        .lut({
            `INST_NUM_WIDTH'd`lui,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`auipc,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`jal,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`jalr,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`beq,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`bne,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`blt,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`bge,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`bltu,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`bgeu,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`lb,
            alu_result,
            `INST_NUM_WIDTH'd`lh,
            alu_result,
            `INST_NUM_WIDTH'd`lw,
            alu_result,
            `INST_NUM_WIDTH'd`lbu,
            alu_result,
            `INST_NUM_WIDTH'd`lhu,
            alu_result,
            `INST_NUM_WIDTH'd`sb,
            alu_result,
            `INST_NUM_WIDTH'd`sh,
            alu_result,
            `INST_NUM_WIDTH'd`sw,
            alu_result,
            `INST_NUM_WIDTH'd`addi,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`slti,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`sltiu,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`xori,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`ori,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`andi,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`slli,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`srli,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`srai,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`add,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`sub,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`sll,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`slt,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`sltu,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`ixor,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`srl,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`sra,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`ior,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`iand,
            `BASE_ADDR,
            `INST_NUM_WIDTH'd`ebreak,
            `BASE_ADDR
        })
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(`MEM_MASK_WIDTH)
    ) muxkeywithdefault_mem_mask (
        .out(mem_mask),
        .key(inst_num),
        .default_out(`MEM_MASK_WIDTH'b0),
        .lut({
            `INST_NUM_WIDTH'd`lui,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`auipc,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`jal,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`jalr,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`beq,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`bne,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`blt,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`bge,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`bltu,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`bgeu,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`lb,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`lh,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`lw,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`lbu,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`lhu,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`sb,
            `MEM_MASK_WIDTH'b0001,
            `INST_NUM_WIDTH'd`sh,
            `MEM_MASK_WIDTH'b0011,
            `INST_NUM_WIDTH'd`sw,
            `MEM_MASK_WIDTH'b1111,
            `INST_NUM_WIDTH'd`addi,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`slti,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`sltiu,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`xori,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`ori,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`andi,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`slli,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`srli,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`srai,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`add,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`sub,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`sll,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`slt,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`sltu,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`ixor,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`srl,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`sra,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`ior,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`iand,
            `MEM_MASK_WIDTH'b0,
            `INST_NUM_WIDTH'd`ebreak,
            `MEM_MASK_WIDTH'b0
        })
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(1)
    ) muxkeywithdefault_mem_r_en (
        .out(mem_r_en),
        .key(inst_num),
        .default_out(1'b0),
        .lut({
            `INST_NUM_WIDTH'd`lui,
            1'b0,
            `INST_NUM_WIDTH'd`auipc,
            1'b0,
            `INST_NUM_WIDTH'd`jal,
            1'b0,
            `INST_NUM_WIDTH'd`jalr,
            1'b0,
            `INST_NUM_WIDTH'd`beq,
            1'b0,
            `INST_NUM_WIDTH'd`bne,
            1'b0,
            `INST_NUM_WIDTH'd`blt,
            1'b0,
            `INST_NUM_WIDTH'd`bge,
            1'b0,
            `INST_NUM_WIDTH'd`bltu,
            1'b0,
            `INST_NUM_WIDTH'd`bgeu,
            1'b0,
            `INST_NUM_WIDTH'd`lb,
            1'b1,
            `INST_NUM_WIDTH'd`lh,
            1'b1,
            `INST_NUM_WIDTH'd`lw,
            1'b1,
            `INST_NUM_WIDTH'd`lbu,
            1'b1,
            `INST_NUM_WIDTH'd`lhu,
            1'b1,
            `INST_NUM_WIDTH'd`sb,
            1'b0,
            `INST_NUM_WIDTH'd`sh,
            1'b0,
            `INST_NUM_WIDTH'd`sw,
            1'b0,
            `INST_NUM_WIDTH'd`addi,
            1'b0,
            `INST_NUM_WIDTH'd`slti,
            1'b0,
            `INST_NUM_WIDTH'd`sltiu,
            1'b0,
            `INST_NUM_WIDTH'd`xori,
            1'b0,
            `INST_NUM_WIDTH'd`ori,
            1'b0,
            `INST_NUM_WIDTH'd`andi,
            1'b0,
            `INST_NUM_WIDTH'd`slli,
            1'b0,
            `INST_NUM_WIDTH'd`srli,
            1'b0,
            `INST_NUM_WIDTH'd`srai,
            1'b0,
            `INST_NUM_WIDTH'd`add,
            1'b0,
            `INST_NUM_WIDTH'd`sub,
            1'b0,
            `INST_NUM_WIDTH'd`sll,
            1'b0,
            `INST_NUM_WIDTH'd`slt,
            1'b0,
            `INST_NUM_WIDTH'd`sltu,
            1'b0,
            `INST_NUM_WIDTH'd`ixor,
            1'b0,
            `INST_NUM_WIDTH'd`srl,
            1'b0,
            `INST_NUM_WIDTH'd`sra,
            1'b0,
            `INST_NUM_WIDTH'd`ior,
            1'b0,
            `INST_NUM_WIDTH'd`iand,
            1'b0,
            `INST_NUM_WIDTH'd`ebreak,
            1'b0
        })
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_TYPE_MAX),
        .KEY_LEN (`INST_TYPE_WIDTH),
        .DATA_LEN(1)
    ) muxkeywithdefault_mem_w_en (
        .out(mem_w_en),
        .key(inst_type),
        .default_out(1'b0),
        .lut({
            `INST_TYPE_WIDTH'd`R,
            1'b0,
            `INST_TYPE_WIDTH'd`I,
            1'b0,
            `INST_TYPE_WIDTH'd`S,
            1'b1,
            `INST_TYPE_WIDTH'd`B,
            1'b0,
            `INST_TYPE_WIDTH'd`U,
            1'b0,
            `INST_TYPE_WIDTH'd`J,
            1'b0
        })
    );

endmodule
