`include "config.vh"
`include "inst.vh"

module exu_alu
    (
        input wire clk,
        input wire rst,
        input wire [`INST_NUM_WIDTH-1:0] inst_num,
        input wire [`INST_TYPE_WIDTH-1:0] inst_type,
        input wire [`IMM_WIDTH-1:0] imm,
        input wire [`SHAMT_WIDTH-1:0] shamt,
        input wire [`ISA_WIDTH-1:0] pc_out,
        input wire [`ISA_WIDTH-1:0] src1,
        input wire [`ISA_WIDTH-1:0] src2,
        input wire [`ISA_WIDTH-1:0] mem_r,
        input wire [`ISA_WIDTH-1:0] alu_result,
        output wire [`ISA_WIDTH-1:0] alu_a,
        output wire [`ISA_WIDTH-1:0] alu_b,
        output wire [`ALU_FUNCT_WIDTH-1:0] alu_funct
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(`ISA_WIDTH)
    ) muxkeywithdefault_alu_a (
        .out(alu_a),
        .key(inst_num),
        .default_out(`ISA_WIDTH'b0),
        .lut({
            `INST_NUM_WIDTH'd`lui,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`auipc,
            pc_out,
            `INST_NUM_WIDTH'd`jal,
            pc_out,
            `INST_NUM_WIDTH'd`jalr,
            pc_out,
            `INST_NUM_WIDTH'd`beq,
            src1,
            `INST_NUM_WIDTH'd`bne,
            src1,
            `INST_NUM_WIDTH'd`bge,
            src1,
            `INST_NUM_WIDTH'd`lw,
            src1,
            `INST_NUM_WIDTH'd`lbu,
            src1,
            `INST_NUM_WIDTH'd`sb,
            src1,
            `INST_NUM_WIDTH'd`sh,
            src1,
            `INST_NUM_WIDTH'd`sw,
            src1,
            `INST_NUM_WIDTH'd`addi,
            src1,
            `INST_NUM_WIDTH'd`sltiu,
            src1,
            `INST_NUM_WIDTH'd`xori,
            src1,
            `INST_NUM_WIDTH'd`andi,
            src1,
            `INST_NUM_WIDTH'd`srai,
            src1,
            `INST_NUM_WIDTH'd`add,
            src1,
            `INST_NUM_WIDTH'd`sub,
            src1,
            `INST_NUM_WIDTH'd`sll,
            src1,
            `INST_NUM_WIDTH'd`sltu,
            src1,
            `INST_NUM_WIDTH'd`ixor,
            src1,
            `INST_NUM_WIDTH'd`ior,
            src1,
            `INST_NUM_WIDTH'd`iand,
            src1,
            `INST_NUM_WIDTH'd`ebreak,
            `ISA_WIDTH'b0
        })
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(`ISA_WIDTH)
    ) muxkeywithdefault_alu_b (
        .out(alu_b),
        .key(inst_num),
        .default_out(`ISA_WIDTH'b0),
        .lut({
            `INST_NUM_WIDTH'd`lui,
            `ISA_WIDTH'b0,
            `INST_NUM_WIDTH'd`auipc,
            imm,
            `INST_NUM_WIDTH'd`jal,
            `ISA_WIDTH'd4,
            `INST_NUM_WIDTH'd`jalr,
            `ISA_WIDTH'd4,
            `INST_NUM_WIDTH'd`beq,
            src2,
            `INST_NUM_WIDTH'd`bne,
            src2,
            `INST_NUM_WIDTH'd`bge,
            src2,
            `INST_NUM_WIDTH'd`lw,
            imm,
            `INST_NUM_WIDTH'd`lbu,
            imm,
            `INST_NUM_WIDTH'd`sb,
            imm,
            `INST_NUM_WIDTH'd`sh,
            imm,
            `INST_NUM_WIDTH'd`sw,
            imm,
            `INST_NUM_WIDTH'd`addi,
            imm,
            `INST_NUM_WIDTH'd`sltiu,
            imm,
            `INST_NUM_WIDTH'd`xori,
            imm,
            `INST_NUM_WIDTH'd`andi,
            imm,
            `INST_NUM_WIDTH'd`srai,
            {{`ISA_WIDTH-`SHAMT_WIDTH{1'b0}},shamt},
            `INST_NUM_WIDTH'd`add,
            src2,
            `INST_NUM_WIDTH'd`sub,
            src2,
            `INST_NUM_WIDTH'd`sll,
            src2,
            `INST_NUM_WIDTH'd`sltu,
            src2,
            `INST_NUM_WIDTH'd`ixor,
            src2,
            `INST_NUM_WIDTH'd`ior,
            src2,
            `INST_NUM_WIDTH'd`iand,
            src2,
            `INST_NUM_WIDTH'd`ebreak,
            `ISA_WIDTH'b0
        })
    );

    MuxKeyWithDefault #(
        .NR_KEY  (`INST_NUM_MAX),
        .KEY_LEN (`INST_NUM_WIDTH),
        .DATA_LEN(`ALU_FUNCT_WIDTH)
    ) muxkeywithdefault_alu_funct (
        .out(alu_funct),
        .key(inst_num),
        .default_out(`ALU_FUNCT_WIDTH'd`NO_FUNCT),
        .lut({
            `INST_NUM_WIDTH'd`auipc,
            `ALU_FUNCT_WIDTH'd`NO_FUNCT,
            `INST_NUM_WIDTH'd`auipc,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`jal,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`jalr,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`beq,
            `ALU_FUNCT_WIDTH'd`EQ,
            `INST_NUM_WIDTH'd`bne,
            `ALU_FUNCT_WIDTH'd`NEQ,
            `INST_NUM_WIDTH'd`bge,
            `ALU_FUNCT_WIDTH'd`GREATER_EQ,
            `INST_NUM_WIDTH'd`lw,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`lbu,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`sb,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`sh,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`sw,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`addi,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`sltiu,
            `ALU_FUNCT_WIDTH'd`LESS_U,
            `INST_NUM_WIDTH'd`xori,
            `ALU_FUNCT_WIDTH'd`XOR,
            `INST_NUM_WIDTH'd`andi,
            `ALU_FUNCT_WIDTH'd`AND,
            `INST_NUM_WIDTH'd`srai,
            `ALU_FUNCT_WIDTH'd`SHIFT_R_A,
            `INST_NUM_WIDTH'd`add,
            `ALU_FUNCT_WIDTH'd`ADD,
            `INST_NUM_WIDTH'd`sub,
            `ALU_FUNCT_WIDTH'd`SUB,
            `INST_NUM_WIDTH'd`sll,
            `ALU_FUNCT_WIDTH'd`SHIFT_L_L,
            `INST_NUM_WIDTH'd`sltu,
            `ALU_FUNCT_WIDTH'd`LESS_U,
            `INST_NUM_WIDTH'd`ixor,
            `ALU_FUNCT_WIDTH'd`XOR,
            `INST_NUM_WIDTH'd`ior,
            `ALU_FUNCT_WIDTH'd`OR,
            `INST_NUM_WIDTH'd`iand,
            `ALU_FUNCT_WIDTH'd`AND,
            `INST_NUM_WIDTH'd`ebreak,
            `ALU_FUNCT_WIDTH'd`NO_FUNCT
        })
    );

endmodule
