`define ysyx_23060075_ISA_WIDTH 32
`define ysyx_23060075_REG_ADDR_WIDTH 4
`define ysyx_23060075_OPCODE_WIDTH 7
`define ysyx_23060075_IMM_WIDTH `ysyx_23060075_ISA_WIDTH
`define ysyx_23060075_SHAMT_WIDTH 5
`define ysyx_23060075_FUNCT3_WIDTH 3
`define ysyx_23060075_FUNCT7_WIDTH 7

`define ysyx_23060075_BASE_ADDR `ysyx_23060075_ISA_WIDTH'h80000000
`define ysyx_23060075_PC_BASE_ADDR `ysyx_23060075_BASE_ADDR
`define ysyx_23060075_MEM_MASK_WIDTH 4

`define ysyx_23060075_ALU_FUNCT_WIDTH 4
`define ysyx_23060075_ALU_FUNCT_MAX 14
`define ysyx_23060075_NO_FUNCT 2
`define ysyx_23060075_ADD 0
`define ysyx_23060075_SUB 8
`define ysyx_23060075_LT 10
`define ysyx_23060075_LTU 11
`define ysyx_23060075_SLL 1
`define ysyx_23060075_SRL 5
`define ysyx_23060075_SRA 13
`define ysyx_23060075_XOR 4
`define ysyx_23060075_OR 6
`define ysyx_23060075_AND 7
`define ysyx_23060075_EQ 9
`define ysyx_23060075_NE 12
`define ysyx_23060075_GE 14
`define ysyx_23060075_GEU 15

`define ysyx_23060075_INST_TYPE_WIDTH 3
`define ysyx_23060075_INST_TYPE_MAX 6
`define ysyx_23060075_N 0
`define ysyx_23060075_R 1
`define ysyx_23060075_I 2
`define ysyx_23060075_S 3
`define ysyx_23060075_B 4
`define ysyx_23060075_U 5
`define ysyx_23060075_J 6

`define ysyx_23060075_OPCODE_NUMBER_MAX 10
