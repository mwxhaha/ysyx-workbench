`define ysyx_23060075_ISA_WIDTH 32
`define ysyx_23060075_IMM_WIDTH `ysyx_23060075_ISA_WIDTH
`define ysyx_23060075_SHAMT_WIDTH 5
`define ysyx_23060075_FUNCT3_WIDTH 3
`define ysyx_23060075_FUNCT7_WIDTH 7

`define ysyx_23060075_BASE_ADDR `ysyx_23060075_ISA_WIDTH'h80000000
`define ysyx_23060075_PC_BASE_ADDR `ysyx_23060075_BASE_ADDR
`define ysyx_23060075_MEM_MASK_WIDTH 4

`define ysyx_23060075_REG_ADDR_WIDTH 4

`define ysyx_23060075_CSR_ADDR_WIDTH 12
`define ysyx_23060075_CSR_ADDR_MEPC `ysyx_23060075_CSR_ADDR_WIDTH'h341
`define ysyx_23060075_CSR_ADDR_MCAUSE `ysyx_23060075_CSR_ADDR_WIDTH'h342
`define ysyx_23060075_CSR_ADDR_MTVEC `ysyx_23060075_CSR_ADDR_WIDTH'h305
`define ysyx_23060075_CSR_ADDR_MSTATUS `ysyx_23060075_CSR_ADDR_WIDTH'h300
`define ysyx_23060075_INTR_CODE_MECALL `ysyx_23060075_ISA_WIDTH'd11
`define ysyx_23060075_MSTATUS_INIT `ysyx_23060075_ISA_WIDTH'h00001800

`define ysyx_23060075_OPCODE_WIDTH 7
`define ysyx_23060075_OPCODE_NUMBER_MAX 10

`define ysyx_23060075_INST_TYPE_WIDTH 3
`define ysyx_23060075_N `ysyx_23060075_INST_TYPE_WIDTH'd0
`define ysyx_23060075_R `ysyx_23060075_INST_TYPE_WIDTH'd1
`define ysyx_23060075_I `ysyx_23060075_INST_TYPE_WIDTH'd2
`define ysyx_23060075_S `ysyx_23060075_INST_TYPE_WIDTH'd3
`define ysyx_23060075_B `ysyx_23060075_INST_TYPE_WIDTH'd4
`define ysyx_23060075_U `ysyx_23060075_INST_TYPE_WIDTH'd5
`define ysyx_23060075_J `ysyx_23060075_INST_TYPE_WIDTH'd6

`define ysyx_23060075_DNPC_MUX_SEL_WIDTH 3
`define ysyx_23060075_DNPC_IS_NO_FUNCT `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b000
`define ysyx_23060075_DNPC_IS_SNPC `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b001
`define ysyx_23060075_DNPC_IS_PC_IMM `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b010
`define ysyx_23060075_DNPC_IS_ALU_RESULT `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b011
`define ysyx_23060075_DNPC_IS_BRANCH `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b100
`define ysyx_23060075_DNPC_IS_MTVEC `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b101
`define ysyx_23060075_DNPC_IS_MEPC `ysyx_23060075_DNPC_MUX_SEL_WIDTH'b110

`define ysyx_23060075_ALU_FUNCT_WIDTH 4
`define ysyx_23060075_NO_FUNCT `ysyx_23060075_ALU_FUNCT_WIDTH'b0010
`define ysyx_23060075_ADD `ysyx_23060075_ALU_FUNCT_WIDTH'b0000
`define ysyx_23060075_SUB `ysyx_23060075_ALU_FUNCT_WIDTH'b1000
`define ysyx_23060075_LT `ysyx_23060075_ALU_FUNCT_WIDTH'b1010
`define ysyx_23060075_LTU `ysyx_23060075_ALU_FUNCT_WIDTH'b1011
`define ysyx_23060075_XOR `ysyx_23060075_ALU_FUNCT_WIDTH'b0100
`define ysyx_23060075_OR `ysyx_23060075_ALU_FUNCT_WIDTH'b0110
`define ysyx_23060075_AND `ysyx_23060075_ALU_FUNCT_WIDTH'b0111
`define ysyx_23060075_SLL `ysyx_23060075_ALU_FUNCT_WIDTH'b0001
`define ysyx_23060075_SRL `ysyx_23060075_ALU_FUNCT_WIDTH'b0101
`define ysyx_23060075_SRA `ysyx_23060075_ALU_FUNCT_WIDTH'b1101
`define ysyx_23060075_EQ `ysyx_23060075_ALU_FUNCT_WIDTH'b1001
`define ysyx_23060075_NE `ysyx_23060075_ALU_FUNCT_WIDTH'b1100
`define ysyx_23060075_GE `ysyx_23060075_ALU_FUNCT_WIDTH'b1110
`define ysyx_23060075_GEU `ysyx_23060075_ALU_FUNCT_WIDTH'b1111

`define ysyx_23060075_SRD_MUX_SEL_WIDTH 3
`define ysyx_23060075_SRD_IS_NO_FUNCT `ysyx_23060075_SRD_MUX_SEL_WIDTH'b000
`define ysyx_23060075_SRD_IS_IMM `ysyx_23060075_SRD_MUX_SEL_WIDTH'b001
`define ysyx_23060075_SRD_IS_PC_IMM `ysyx_23060075_SRD_MUX_SEL_WIDTH'b010
`define ysyx_23060075_SRD_IS_SNPC `ysyx_23060075_SRD_MUX_SEL_WIDTH'b011
`define ysyx_23060075_SRD_IS_MEM_R `ysyx_23060075_SRD_MUX_SEL_WIDTH'b100
`define ysyx_23060075_SRD_IS_ALU_RESULT `ysyx_23060075_SRD_MUX_SEL_WIDTH'b101
`define ysyx_23060075_SRD_IS_CSR_R `ysyx_23060075_SRD_MUX_SEL_WIDTH'b110

`define ysyx_23060075_AXI_MTOS_WIDTH `ysyx_23060075_ISA_WIDTH*3+`ysyx_23060075_MEM_MASK_WIDTH+5
`define ysyx_23060075_AXI_STOM_WIDTH `ysyx_23060075_ISA_WIDTH*3+5
